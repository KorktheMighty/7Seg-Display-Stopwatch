----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/22/2021 02:13:30 AM
-- Design Name: 
-- Module Name: modecontrol - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity modecontrol is
  Port (
        clk,reset,st : in STD_LOGIC;
        
        en           : out STD_LOGIC );
end modecontrol;



architecture Behavioral of modecontrol is

signal mode : STD_LOGIC ;
signal lst  : STD_LOGIC ;
begin
en <= mode;
  process (clk, reset) begin
    if (reset = '1') then
      mode <= '0';
    elsif rising_edge(clk) then
      if (st = '1') and (lst = '0') then
        mode <= not mode;
      end if;
      lst <= st;
    end if;
  end process;


end Behavioral;
